--@ Copyright (c) 2020 Bluespec, Inc. All rights reserved.
--@ 
--@ Redistribution and use in source and binary forms, with or without
--@ modification, are permitted provided that the following conditions are
--@ met:
--@ 
--@ 1. Redistributions of source code must retain the above copyright
--@    notice, this list of conditions and the following disclaimer.
--@ 
--@ 2. Redistributions in binary form must reproduce the above copyright
--@    notice, this list of conditions and the following disclaimer in the
--@    documentation and/or other materials provided with the
--@    distribution.
--@ 
--@ 3. Neither the name of the copyright holder nor the names of its
--@    contributors may be used to endorse or promote products derived
--@    from this software without specific prior written permission.
--@ 
--@ THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
--@ "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
--@ LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
--@ A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT
--@ HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
--@ SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
--@ LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
--@ DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
--@ THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
--@ (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
--@ OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

package ClientServerS(
        ClientS(..), ServerS(..), ClientServerS(..), mkRequestResponseBufferS,
        mkSizedRequestResponseBufferS, mkResponseBufferS, mkRequestBufferS,
        mkRequestResponseBufferS1S, joinServerSsBC, joinServerSs, splitServerS,
        fifosToServerS, fifosToClientS, fifosToClientServerS,
        toGPClientS, toGPServerS)
    where
import qualified Vector
import List
import FIFO
import Counter
import Connectable
import GetPut
import Clocks

--@ \subsubsection{ClientServerS}
--@ \index{ClientServerS@\te{ClientServerS} (package)|textbf}
--@
--@ The interfaces \te{ClientS} and \te{ServerS} can be used for
--@ modules that have a request-response type of interface
--@ (e.g. a RAM).
--@ The ServerS accepts requests and generates responses, and
--@ vice versa for the ClientS.
--@ There are no assumptions about how many (if any) responses
--@ a request will generate.

--@ \index{ClientS@\te{ClientS} (interface)|textbf}
--@ \begin{libverbatim}
--@ interface ClientS #(type a, type b);
--@     interface Get#(a) request();
--@     interface Put#(b) response();
--@ endinterface: ClientS
--@ \end{libverbatim}
interface ClientS a b =
    request  :: Get a
    response :: Put b

--@ \index{ServerS@\te{ServerS} (interface)|textbf}
--@ \begin{libverbatim}
--@ interface ServerS #(type a, type b);
--@     interface Put#(a) request();
--@     interface Get#(b) response();
--@ endinterface: ServerS
--@ \end{libverbatim}
interface ServerS a b =
    request  :: Put a
    response :: Get b

--@ A \te{ClientS} can be connected to a \te{ServerS}
--@ and vice versa.
--@ \begin{libverbatim}
--@ instance Connectable #(ClientS#(a, b), ServerS#(a, b));
--@ instance Connectable #(ServerS#(a, b), ClientS#(a, b));
--@ \end{libverbatim}
instance Connectable (ClientS a b) (ServerS a b)
   where
    mkConnection :: (IsModule m c ) => ClientS a b -> ServerS a b -> m Empty
    mkConnection c s =
       module
          rules
            "ClientServerSRequest":when True
             ==> action
                    x :: a <- c.request.get
                    s.request.put x
            "ClientServerSResponse":when True
             ==> action
                    x :: b <- s.response.get
                    c.response.put x

instance Connectable (ServerS a b) (ClientS a b)
   where
    mkConnection s c = mkConnection c s

instance (Bits a sa, Bits b sb) => ClockConv (ClientS a b) where
    mkConverter :: (Prelude.IsModule m c) => Integer -> ClientS a b -> m (ClientS a b)
    mkConverter d cluses =
        module
            req  <- mkConverter d cluses.request
            resp <- mkConverter d cluses.response

            interface
              request  = req
              response = resp

instance (Bits a sa, Bits b sb) => ClockConv (ServerS a b) where
    mkConverter :: (Prelude.IsModule m c) => Integer -> ServerS a b -> m (ServerS a b)
    mkConverter d cluses =
        module
            req  <- mkConverter d cluses.request
            resp <- mkConverter d cluses.response

            interface
              request  = req
              response = resp

--@ \lineup
--@ \begin{libverbatim}
--@ typedef Tuple2 #(ClientS#(a, b), ServerS#(a, b)) ClientServerS #(type a, type b);
--@ \end{libverbatim}
type ClientServerS a b = (ClientS a b, ServerS a b)

--@ Create a buffer that just passes requests and responses between the
--@ two generated interfaces.
--@ \index{mkRequestResponseBufferS@\te{mkRequestResponseBufferS} (function)|textbf}
--@ \begin{libverbatim}
--@ module mkRequestResponseBufferS(ClientServerS#(a, b))
--@   provisos (Bits#(a, sa), Bits#(b, sb));
--@ \end{libverbatim}
mkRequestResponseBufferS :: (IsModule m c , Bits a sa, Bits b sb) => m (ClientServerS a b)
mkRequestResponseBufferS =
    module
        (qget, qput) :: (Get a, Put a) <- mkGetPut
        (sget, sput) :: (Get b, Put b) <- mkGetPut
        let c = interface ClientS
                    request  = qget
                    response = sput
            s = interface ServerS
                    request  = qput
                    response = sget
        interface (c, s)

--@ Create a buffer that just passes requests and responses between the
--@ two generated interfaces.  Uses half the flops of
--@ \te{mkRequestResponseBufferS}, but also has half the throughput.
--@ \index{mkRequestResponseBufferS1S@\te{mkRequestResponseBufferS1S} (function)|textbf}
--@ \begin{libverbatim}
--@ module mkRequestResponseBufferS1S(ClientServerS#(a, b))
--@   provisos (Bits#(a, sa), Bits#(b, sb));
--@ \end{libverbatim}
mkRequestResponseBufferS1S :: (IsModule m c , Bits a sa, Bits b sb) => m (ClientServerS a b)
mkRequestResponseBufferS1S =
    module
        (qget, qput) :: (Get a, Put a) <- mkGPFIFO1
        (sget, sput) :: (Get b, Put b) <- mkGPFIFO1
        let c = interface ClientS
                    request  = qget
                    response = sput
            s = interface ServerS
                    request  = qput
                    response = sget
        interface (c, s)

--@ The same, using sized FIFOs.
--@ \index{mkSizedRequestResponseBufferS@\te{mkSizedRequestResponseBufferS} (function)|textbf}
--@ \begin{libverbatim}
--@ module mkSizedRequestResponseBufferS#(Integer sz)(ClientServerS#(a, b))
--@   provisos (Bits#(a, sa), Bits#(b, sb));
--@ \end{libverbatim}
mkSizedRequestResponseBufferS :: (IsModule m c , Bits a sa, Bits b sb) => Integer -> m (ClientServerS a b)
mkSizedRequestResponseBufferS sz =
    module
        (qget, qput) :: (Get a, Put a) <- mkGPSizedFIFO sz
        (sget, sput) :: (Get b, Put b) <- mkGPSizedFIFO sz
        let c = interface ClientS
                    request  = qget
                    response = sput
            s = interface ServerS
                    request  = qput
                    response = sget
        interface (c, s)


--@ Create a new ServerS with buffered requests.
--@ \index{mkRequestBufferS@\te{mkRequestBufferS} (function)|textbf}
--@ \begin{libverbatim}
--@ module mkRequestBufferS#(ServerS#(a, b) s)(ServerS#(a, b))
--@   provisos (Bits#(a, sa));
--@ \end{libverbatim}
mkRequestBufferS :: (IsModule m c , Bits a sa) => ServerS a b -> m (ServerS a b)
mkRequestBufferS s =
    module
        (qget, qput) :: (Get a, Put a) <- mkGetPut
        rules
              "mkRequestBufferS" : when True ==>
                 action
                   x :: a <- qget.get
                   s.request.put x

        interface -- ServerS
                    request  = qput
                    response = s.response


--@ Create a new ServerS with buffered responses.
--@ \index{mkResponseBufferS@\te{mkResponseBufferS} (function)|textbf}
--@ \begin{libverbatim}
--@ module mkResponseBufferS#(ServerS#(a, b) s)(ServerS#(a, b))
--@   provisos (Bits#(b, sb));
--@ \end{libverbatim}
mkResponseBufferS :: (IsModule m c , Bits b sb) => ServerS a b -> m (ServerS a b)
mkResponseBufferS s =
    module
        (sget, sput) :: (Get b, Put b) <- mkGetPut
        rules
              "mkResponseBufferS" : when True ==>
                 action
                   x :: b <- s.response.get
                   sput.put x

        interface -- ServerS
                    request  = s.request
                    response = sget

--@ Join a list of ServerS's to one ServerS.  All incoming requests are broadcasted
--@ all the ServerS's and all responses are merged.
--@ The function introduces a one cycle latency on the response.
--@ \index{joinServerSsSBC@\te{joinServerSsSBC} (function)|textbf}
--@ \begin{libverbatim}
--@ module joinServerSsSBC#(List#(ServerS#(a, b)) ifs)(ServerS#(a, b))
--@   provisos (Bits#(b, sb));
--@ \end{libverbatim}
joinServerSsBC :: (IsModule m c , Bits b sb) => List (ServerS a b) -> m (ServerS a b)
joinServerSsBC ifs =
  module
    (sget, sput) :: (Get b, Put b) <- mkGetPut
    let rl s =
            rules
              "joinServerSsSBC":
                when True ==>
                 action
                   x <- (s :: ServerS a b).response.get
                   sput.put x
    addRules $ foldr (<+>) (rules {}) (map rl ifs)
    interface -- ServerS
            request =
             interface Put
              put req = joinActions (map (\ i -> (i :: ServerS a b).request.put req) ifs)
            response = sget

--@ Join a list of ServerSs to one ServerS.  All incoming requests are sent to
--@ a selected subset of the ServerSs and all responses are merged.
--@ The selection is my a function that can transform the request type
--@ while testing if it should be sent on.
--@ The function introduces a one cycle latency on the response.
--@ \index{joinServerSs@\te{joinServerSs} (function)|textbf}
--@ \begin{libverbatim}
--@ module joinServerSs#( List#(Tuple2 #(a -> Maybe#(a'),
--@                      ServerS#(a', b))) ifs)(ServerS#(a, b))
--@   provisos (Bits#(b, sb));
--@ \end{libverbatim}
joinServerSs ::  (IsModule m c , Bits b sb) => List (a -> Maybe a', ServerS a' b) -> m (ServerS a b)
joinServerSs ifs =
  module
    (sget, sput) :: (Get b, Put b) <- mkGetPut
    let rl (_, s) =
            rules
              "joinServerSs":
                when True ==>
                  action
                   x <- (s :: ServerS a' b).response.get
                   sput.put x
        send req (f, s) =
            case f req of
            Nothing -> noAction
            Just req' -> (s :: ServerS a' b).request.put req'
    addRules $ foldr (<+>) (rules {}) (map rl ifs)
    interface -- ServerS
            request =
             interface Put
              put req = joinActions (map (send req) ifs)
            response = sget

type MaxLat = 8        -- XXX This is just wrong
--@ Split a ServerS into a number of identical ServerSs.
--@ The integer argument specifies how many outstanding requests
--@ a returned ServerS may have.  This number should be
--@ the latency of the argument ServerS to sustain full bandwidth.
--@ (A small number still works, as does a larger number.)
--@ \index{splitServerS@\te{splitServerS} (function)|textbf}
--@ \begin{libverbatim}
--@ module splitServerS#(Integer lat, ServerS#(a, b) serv)(Vector#(n, ServerS#(a, b)))
--@   provisos (Bits#(b, sb), Log#(n, ln));
--@ \end{libverbatim}
splitServerS :: (IsModule m c , Bits b sb, Log n ln) =>
               Integer -> ServerS a b -> m (Vector.Vector n (ServerS a b))
splitServerS lat serv =
  module
    tags :: FIFO (Bit ln) <- mkSizedFIFO lat
    let mkServ :: (Bit ln) -> m (ServerS a b)
        mkServ i =
          module
            out :: FIFO b <- mkSizedFIFO lat
            cnt :: Counter MaxLat <- mkCounter (fromInteger lat)
            rules
                when tags.first == i
                 ==> action
                        tags.deq
                        x <- serv.response.get
                        out.enq x
            interface ServerS
              request =
                interface Put
                  put req =
                        action
                            serv.request.put req
                            tags.enq i
                            cnt.down
                    when cnt.value > 0
              response =
                interface Get
                  get = do
                            out.deq
                            cnt.up
                            return out.first
    Vector.mapM (mkServ ∘ fromInteger) Vector.genList

--@ fifosToServerS

fifosToServerS :: FIFO rq -> FIFO rs -> ServerS rq rs
fifosToServerS rqf rsf =
    interface ServerS
       request  = fifoToPut rqf
       response = fifoToGet rsf

fifosToClientS :: FIFO rq -> FIFO rs -> ClientS rq rs
fifosToClientS rqf rsf =
    interface ClientS
       request  = fifoToGet rqf
       response = fifoToPut rsf

fifosToClientServerS :: FIFO rq -> FIFO rs -> ClientServerS rq rs
fifosToClientServerS rqf rsf = (fifosToClientS rqf rsf, fifosToServerS rqf rsf)

-- toGPClientS, toGPServerS

toGPClientS :: (ToGet rq_ifc rq, ToPut rs_ifc rs) =>
              rq_ifc -> rs_ifc -> ClientS rq rs
toGPClientS rqi rsi =
    interface ClientS
        request = toGet rqi
        response = toPut rsi

toGPServerS :: (ToPut rq_ifc rq, ToGet rs_ifc rs) =>
              rq_ifc -> rs_ifc -> ServerS rq rs
toGPServerS rqi rsi =
    interface ServerS
        request = toPut rqi
        response = toGet rsi

