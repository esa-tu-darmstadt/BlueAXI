package BlueAXI;

import AXI4_Lite :: *;
import GenericAxi4LiteSlave :: *;

import AXI4 :: *;
import AXI4_Stream :: *;
import GenericAxi4Master :: *;

import BlueAXITests :: *;
import BlueAXIBRAM :: *;

import AXI4_Monitor :: *;

import AXI3 :: *;

export AXI4_Lite :: *;
export GenericAxi4LiteSlave :: *;

export AXI4 :: *;
export GenericAxi4Master :: *;

export BlueAXITests :: *;
export BlueAXIBRAM :: *;

export AXI4_Monitor :: *;

export AXI3 :: *;

endpackage